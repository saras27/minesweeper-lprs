
-------------------------------------------------------
-- Logicko projektovanje racunarskih sistema 1
-- 2011/2012,2020
--
-- Instruction ROM
--
-- author:
-- Ivan Kastelan (ivan.kastelan@rt-rk.com)
-- Milos Subotic (milos.subotic@uns.ac.rs)
-------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity instr_rom is
	port(
		iA : in  std_logic_vector(15 downto 0);
		oQ : out std_logic_vector(14 downto 0)
	);
end entity instr_rom;

-- ubaciti sadrzaj *.txt datoteke generisane pomocu lprsasm ------
architecture Behavioral of instr_rom is
begin
    oQ <= "000010000000000"  when iA = 0 else
          "000110000000000"  when iA = 1 else
          "000110000000000"  when iA = 2 else
          "000110000000000"  when iA = 3 else
          "000110000000000"  when iA = 4 else
          "100000111000000"  when iA = 5 else
          "000110000000000"  when iA = 6 else
          "000110000000000"  when iA = 7 else
          "100000101000000"  when iA = 8 else
          "000010000000000"  when iA = 9 else
          "000110001000000"  when iA = 10 else
          "100000000000000"  when iA = 11 else
          "000000011000000"  when iA = 12 else
          "000110000000000"  when iA = 13 else
          "000110000000000"  when iA = 14 else
          "100000001000001"  when iA = 15 else
          "001000001001000"  when iA = 16 else
          "000010001001000"  when iA = 17 else
          "100000001000001"  when iA = 18 else
          "001000110011000"  when iA = 19 else
          "001000110110000"  when iA = 20 else
          "001000110110000"  when iA = 21 else
          "000111110110000"  when iA = 22 else
          "100000010000000"  when iA = 23 else
          "010010000100110"  when iA = 24 else
          "000010100010011"  when iA = 25 else
          "010101000100100"  when iA = 26 else
          "110000000100000"  when iA = 27 else
          "000001100001000"  when iA = 28 else
          "000011100100110"  when iA = 29 else
          "000001100100011"  when iA = 30 else
          "000110100100000"  when iA = 31 else
          "000110100100000"  when iA = 32 else
          "110000000011100"  when iA = 33 else
          "001000001001000"  when iA = 34 else
          "000110001001000"  when iA = 35 else
          "000110000000000"  when iA = 36 else
          "010000000010111"  when iA = 37 else
          "000010000000000"  when iA = 38 else
          "000110000000000"  when iA = 39 else
          "100000000000000"  when iA = 40 else
          "000010010010010"  when iA = 41 else
          "100000001000000"  when iA = 42 else
          "010010000101111"  when iA = 43 else
          "110000000010000"  when iA = 44 else
          "000110000000000"  when iA = 45 else
          "010000000101010"  when iA = 46 else
          "000010000000000"  when iA = 47 else
          "100000000000000"  when iA = 48 else
          "000110000000000"  when iA = 49 else
          "000110000000000"  when iA = 50 else
          "000010011011011"  when iA = 51 else
          "100000011000011"  when iA = 52 else
          "000010001001001"  when iA = 53 else
          "100000010000000"  when iA = 54 else
          "010010000111101"  when iA = 55 else
          "000010100010011"  when iA = 56 else
          "010001000111011"  when iA = 57 else
          "110000000001000"  when iA = 58 else
          "000110000000000"  when iA = 59 else
          "010000000110110"  when iA = 60 else
          "000010000000000"  when iA = 61 else
          "100000000000000"  when iA = 62 else
          "000000001000000"  when iA = 63 else
          "000110000000000"  when iA = 64 else
          "000110000000000"  when iA = 65 else
          "100000010000000"  when iA = 66 else
          "010010010101011"  when iA = 67 else
          "000010011010001"  when iA = 68 else
          "010101010101001"  when iA = 69 else
          "000000100001000"  when iA = 70 else
          "000110100100000"  when iA = 71 else
          "000110100100000"  when iA = 72 else
          "000010100000100"  when iA = 73 else
          "000000010001000"  when iA = 74 else
          "000111010010000"  when iA = 75 else
          "000011010010100"  when iA = 76 else
          "000000011100000"  when iA = 77 else
          "001001011011000"  when iA = 78 else
          "001001011011000"  when iA = 79 else
          "001001011011000"  when iA = 80 else
          "000000011011000"  when iA = 81 else
          "010001001110001"  when iA = 82 else
          "000010000000001"  when iA = 83 else
          "100000100000000"  when iA = 84 else
          "000010100100001"  when iA = 85 else
          "010001001011010"  when iA = 86 else
          "100000100000000"  when iA = 87 else
          "000110100100000"  when iA = 88 else
          "110000000100000"  when iA = 89 else
          "000000010010000"  when iA = 90 else
          "010001001100100"  when iA = 91 else
          "000111000000000"  when iA = 92 else
          "100000100000000"  when iA = 93 else
          "000010100100001"  when iA = 94 else
          "010001001100011"  when iA = 95 else
          "100000100000000"  when iA = 96 else
          "000110100100000"  when iA = 97 else
          "110000000100000"  when iA = 98 else
          "000110000000000"  when iA = 99 else
          "000000100010000"  when iA = 100 else
          "000110100100000"  when iA = 101 else
          "000010100100001"  when iA = 102 else
          "010001001110000"  when iA = 103 else
          "000110000000000"  when iA = 104 else
          "100000100000000"  when iA = 105 else
          "000010100100001"  when iA = 106 else
          "010001001101111"  when iA = 107 else
          "100000100000000"  when iA = 108 else
          "000110100100000"  when iA = 109 else
          "110000000100000"  when iA = 110 else
          "000111000000000"  when iA = 111 else
          "000001000000001"  when iA = 112 else
          "000000010010000"  when iA = 113 else
          "010001001111011"  when iA = 114 else
          "000111000000000"  when iA = 115 else
          "100000100000000"  when iA = 116 else
          "000010100100001"  when iA = 117 else
          "010001001111010"  when iA = 118 else
          "100000100000000"  when iA = 119 else
          "000110100100000"  when iA = 120 else
          "110000000100000"  when iA = 121 else
          "000110000000000"  when iA = 122 else
          "000000100010000"  when iA = 123 else
          "000110100100000"  when iA = 124 else
          "000010100100001"  when iA = 125 else
          "010001010000111"  when iA = 126 else
          "000110000000000"  when iA = 127 else
          "100000100000000"  when iA = 128 else
          "000010100100001"  when iA = 129 else
          "010001010000110"  when iA = 130 else
          "100000100000000"  when iA = 131 else
          "000110100100000"  when iA = 132 else
          "110000000100000"  when iA = 133 else
          "000111000000000"  when iA = 134 else
          "000000100011000"  when iA = 135 else
          "000110100100000"  when iA = 136 else
          "000010100100001"  when iA = 137 else
          "010001010101001"  when iA = 138 else
          "000001000000001"  when iA = 139 else
          "100000100000000"  when iA = 140 else
          "000010100100001"  when iA = 141 else
          "010001010010010"  when iA = 142 else
          "100000100000000"  when iA = 143 else
          "000110100100000"  when iA = 144 else
          "110000000100000"  when iA = 145 else
          "000000010010000"  when iA = 146 else
          "010001010011100"  when iA = 147 else
          "000111000000000"  when iA = 148 else
          "100000100000000"  when iA = 149 else
          "000010100100001"  when iA = 150 else
          "010001010011011"  when iA = 151 else
          "100000100000000"  when iA = 152 else
          "000110100100000"  when iA = 153 else
          "110000000100000"  when iA = 154 else
          "000110000000000"  when iA = 155 else
          "000000100010000"  when iA = 156 else
          "000110100100000"  when iA = 157 else
          "000010100100001"  when iA = 158 else
          "010001010101000"  when iA = 159 else
          "000110000000000"  when iA = 160 else
          "100000100000000"  when iA = 161 else
          "000010100100001"  when iA = 162 else
          "010001010100111"  when iA = 163 else
          "100000100000000"  when iA = 164 else
          "000110100100000"  when iA = 165 else
          "110000000100000"  when iA = 166 else
          "000111000000000"  when iA = 167 else
          "000010000000001"  when iA = 168 else
          "000110000000000"  when iA = 169 else
          "010000001000010"  when iA = 170 else
          "000010110110110"  when iA = 171 else
          "100000110000110"  when iA = 172 else
          "000111110110000"  when iA = 173 else
          "000111110110000"  when iA = 174 else
          "000111110110000"  when iA = 175 else
          "100000110000110"  when iA = 176 else
          "100000000000110"  when iA = 177 else
          "010101010110001"  when iA = 178 else
          "100000000000110"  when iA = 179 else
          "010001010110011"  when iA = 180 else
          "000010011011011"  when iA = 181 else
          "000010000000000"  when iA = 182 else
          "100000000000000"  when iA = 183 else
          "001001111000000"  when iA = 184 else
          "100000111000111"  when iA = 185 else
          "000110000000000"  when iA = 186 else
          "000110000000000"  when iA = 187 else
          "000000001000000"  when iA = 188 else
          "000010100100100"  when iA = 189 else
          "100000100000100"  when iA = 190 else
          "001000100100000"  when iA = 191 else
          "001000100100000"  when iA = 192 else
          "001000100100000"  when iA = 193 else
          "000110100100000"  when iA = 194 else
          "000001011100000"  when iA = 195 else
          "100000011000011"  when iA = 196 else
          "010001011001101"  when iA = 197 else
          "000000011011000"  when iA = 198 else
          "010010011001111"  when iA = 199 else
          "100000011000000"  when iA = 200 else
          "010010011001111"  when iA = 201 else
          "000010010000001"  when iA = 202 else
          "000001010010111"  when iA = 203 else
          "110000000011010"  when iA = 204 else
          "000110000000000"  when iA = 205 else
          "010000011000011"  when iA = 206 else
          "000010111111111"  when iA = 207 else
          "100000111000111"  when iA = 208 else
          "001001111111000"  when iA = 209 else
          "100000111000111"  when iA = 210 else
          "000010000000000"  when iA = 211 else
          "000010011011011"  when iA = 212 else
          "100000011000011"  when iA = 213 else
          "000111011011000"  when iA = 214 else
          "100000000000000"  when iA = 215 else
          "100000001000000"  when iA = 216 else
          "000110000000000"  when iA = 217 else
          "100000010000000"  when iA = 218 else
          "001000010010000"  when iA = 219 else
          "001000010010000"  when iA = 220 else
          "001000010010000"  when iA = 221 else
          "000001010010001"  when iA = 222 else
          "000001010010111"  when iA = 223 else
          "110000000011010"  when iA = 224 else
          "000010000000000"  when iA = 225 else
          "000110000000000"  when iA = 226 else
          "000110000000000"  when iA = 227 else
          "100000001000000"  when iA = 228 else
          "000110000000000"  when iA = 229 else
          "100000010000000"  when iA = 230 else
          "000111000000000"  when iA = 231 else
          "000110001001000"  when iA = 232 else
          "000010010010001"  when iA = 233 else
          "010001011101101"  when iA = 234 else
          "110000000001000"  when iA = 235 else
          "010000010101011"  when iA = 236 else
          "000010001001001"  when iA = 237 else
          "110000000001000"  when iA = 238 else
          "100000000000101"  when iA = 239 else
          "000000000000000"  when iA = 240 else
          "010001110101010"  when iA = 241 else
          "000010000000000"  when iA = 242 else
          "100000000000000"  when iA = 243 else
          "100000001000000"  when iA = 244 else
          "000110000000000"  when iA = 245 else
          "100000010000000"  when iA = 246 else
          "000000100010000"  when iA = 247 else
          "001000100100000"  when iA = 248 else
          "001000100100000"  when iA = 249 else
          "001000100100000"  when iA = 250 else
          "000001100100001"  when iA = 251 else
          "000010000000000"  when iA = 252 else
          "100000000000000"  when iA = 253 else
          "000000011000000"  when iA = 254 else
          "000110011011000"  when iA = 255 else
          "000110011011000"  when iA = 256 else
          "001000000000000"  when iA = 257 else
          "001000000000000"  when iA = 258 else
          "001000000000000"  when iA = 259 else
          "001000000000000"  when iA = 260 else
          "000001000000011"  when iA = 261 else
          "000110000000000"  when iA = 262 else
          "000110000000000"  when iA = 263 else
          "110000000100000"  when iA = 264 else
          "000010000000000"  when iA = 265 else
          "100000000000000"  when iA = 266 else
          "000110000000000"  when iA = 267 else
          "000110000000000"  when iA = 268 else
          "000001100100000"  when iA = 269 else
          "100000000000100"  when iA = 270 else
          "000010001001001"  when iA = 271 else
          "100000001000001"  when iA = 272 else
          "000010001000001"  when iA = 273 else
          "010001111101011"  when iA = 274 else
          "000010000000000"  when iA = 275 else
          "100000000000000"  when iA = 276 else
          "000111000000000"  when iA = 277 else
          "000000011000000"  when iA = 278 else
          "100000000000000"  when iA = 279 else
          "000110000000000"  when iA = 280 else
          "110000000100000"  when iA = 281 else
          "110000000000011"  when iA = 282 else
          "000010000000000"  when iA = 283 else
          "100000000000000"  when iA = 284 else
          "000111000000000"  when iA = 285 else
          "100000001000000"  when iA = 286 else
          "100000010000001"  when iA = 287 else
          "010010110100001"  when iA = 288 else
          "000010000000000"  when iA = 289 else
          "100000000000000"  when iA = 290 else
          "000111000000000"  when iA = 291 else
          "100000001000000"  when iA = 292 else
          "000111001001000"  when iA = 293 else
          "110000000001000"  when iA = 294 else
          "100000011000010"  when iA = 295 else
          "000010100100100"  when iA = 296 else
          "100000100000100"  when iA = 297 else
          "000010100011100"  when iA = 298 else
          "010001110100000"  when iA = 299 else
          "000010001001001"  when iA = 300 else
          "100000001000001"  when iA = 301 else
          "001000001001000"  when iA = 302 else
          "001000001001000"  when iA = 303 else
          "001000001001000"  when iA = 304 else
          "000110001001000"  when iA = 305 else
          "000001001001010"  when iA = 306 else
          "100000100000001"  when iA = 307 else
          "010101110100000"  when iA = 308 else
          "000000011011000"  when iA = 309 else
          "010101110010110"  when iA = 310 else
          "000010000000000"  when iA = 311 else
          "100000000000000"  when iA = 312 else
          "000110000000000"  when iA = 313 else
          "000110000000000"  when iA = 314 else
          "000010000010000"  when iA = 315 else
          "000010011011011"  when iA = 316 else
          "100000011000011"  when iA = 317 else
          "000111011011000"  when iA = 318 else
          "000011011011000"  when iA = 319 else
          "000000100000000"  when iA = 320 else
          "001001100100000"  when iA = 321 else
          "001001100100000"  when iA = 322 else
          "001001100100000"  when iA = 323 else
          "000010110110110"  when iA = 324 else
          "100000110000110"  when iA = 325 else
          "001000110110000"  when iA = 326 else
          "001000110110000"  when iA = 327 else
          "001000110110000"  when iA = 328 else
          "000110110110000"  when iA = 329 else
          "000000100100000"  when iA = 330 else
          "010001101011101"  when iA = 331 else
          "000000000010000"  when iA = 332 else
          "000010001001001"  when iA = 333 else
          "100000001000001"  when iA = 334 else
          "000010000000001"  when iA = 335 else
          "000001001000110"  when iA = 336 else
          "100000001000001"  when iA = 337 else
          "010101101011101"  when iA = 338 else
          "000010001001001"  when iA = 339 else
          "100000001000001"  when iA = 340 else
          "000111001001000"  when iA = 341 else
          "100000001000001"  when iA = 342 else
          "000110001001000"  when iA = 343 else
          "110000000000001"  when iA = 344 else
          "000010000000000"  when iA = 345 else
          "100000000000000"  when iA = 346 else
          "000111000000000"  when iA = 347 else
          "110000000001000"  when iA = 348 else
          "000000011011000"  when iA = 349 else
          "010001101101101"  when iA = 350 else
          "000111000010000"  when iA = 351 else
          "000001001000110"  when iA = 352 else
          "100000001000001"  when iA = 353 else
          "010101101101101"  when iA = 354 else
          "000010001001001"  when iA = 355 else
          "100000001000001"  when iA = 356 else
          "000111001001000"  when iA = 357 else
          "100000001000001"  when iA = 358 else
          "000110001001000"  when iA = 359 else
          "110000000000001"  when iA = 360 else
          "000010000000000"  when iA = 361 else
          "100000000000000"  when iA = 362 else
          "000111000000000"  when iA = 363 else
          "110000000001000"  when iA = 364 else
          "000010001001001"  when iA = 365 else
          "100000001000001"  when iA = 366 else
          "000110000011000"  when iA = 367 else
          "000010000000001"  when iA = 368 else
          "010001110000000"  when iA = 369 else
          "000110000010000"  when iA = 370 else
          "000001001000110"  when iA = 371 else
          "100000001000001"  when iA = 372 else
          "010101110000000"  when iA = 373 else
          "000010001001001"  when iA = 374 else
          "100000001000001"  when iA = 375 else
          "000111001001000"  when iA = 376 else
          "100000001000001"  when iA = 377 else
          "000110001001000"  when iA = 378 else
          "110000000000001"  when iA = 379 else
          "000010000000000"  when iA = 380 else
          "100000000000000"  when iA = 381 else
          "000111000000000"  when iA = 382 else
          "110000000001000"  when iA = 383 else
          "000010000000000"  when iA = 384 else
          "100000000000000"  when iA = 385 else
          "000110001100000"  when iA = 386 else
          "000010000001000"  when iA = 387 else
          "010001110010110"  when iA = 388 else
          "000000000010000"  when iA = 389 else
          "000010001001001"  when iA = 390 else
          "100000001000001"  when iA = 391 else
          "000001000000001"  when iA = 392 else
          "000001001000110"  when iA = 393 else
          "100000001000001"  when iA = 394 else
          "010101110010110"  when iA = 395 else
          "000010001001001"  when iA = 396 else
          "100000001000001"  when iA = 397 else
          "000111001001000"  when iA = 398 else
          "100000001000001"  when iA = 399 else
          "000110001001000"  when iA = 400 else
          "110000000000001"  when iA = 401 else
          "000010000000000"  when iA = 402 else
          "100000000000000"  when iA = 403 else
          "000111000000000"  when iA = 404 else
          "110000000001000"  when iA = 405 else
          "000010001001001"  when iA = 406 else
          "100000001000001"  when iA = 407 else
          "001000001001000"  when iA = 408 else
          "001000001001000"  when iA = 409 else
          "001000001001000"  when iA = 410 else
          "000110001001000"  when iA = 411 else
          "000001001001010"  when iA = 412 else
          "000010100100100"  when iA = 413 else
          "000110100100000"  when iA = 414 else
          "110000000100001"  when iA = 415 else
          "010000100011011"  when iA = 416 else
          "000010000000000"  when iA = 417 else
          "000010001001001"  when iA = 418 else
          "000010001010010"  when iA = 419 else
          "000010001011011"  when iA = 420 else
          "000010100100100"  when iA = 421 else
          "000010111111111"  when iA = 422 else
          "100000111000111"  when iA = 423 else
          "001001111111000"  when iA = 424 else
          "100000111000111"  when iA = 425 else
          "000111101101000"  when iA = 426 else
          "100000010000101"  when iA = 427 else
          "000111101101000"  when iA = 428 else
          "100000001000101"  when iA = 429 else
          "000110101101000"  when iA = 430 else
          "000110101101000"  when iA = 431 else
          "000010000000000"  when iA = 432 else
          "100000000000000"  when iA = 433 else
          "100000011000000"  when iA = 434 else
          "000110000000000"  when iA = 435 else
          "100000100000000"  when iA = 436 else
          "000001011011001"  when iA = 437 else
          "010110110111001"  when iA = 438 else
          "000010011011011"  when iA = 439 else
          "010000111000010"  when iA = 440 else
          "000010000000000"  when iA = 441 else
          "100000000000000"  when iA = 442 else
          "000111000000000"  when iA = 443 else
          "000010000000011"  when iA = 444 else
          "010110111000010"  when iA = 445 else
          "000010011011011"  when iA = 446 else
          "100000011000011"  when iA = 447 else
          "000111011011000"  when iA = 448 else
          "010000111000010"  when iA = 449 else
          "000001100100010"  when iA = 450 else
          "010110111000110"  when iA = 451 else
          "000010100100100"  when iA = 452 else
          "010000111001111"  when iA = 453 else
          "000010000000000"  when iA = 454 else
          "100000000000000"  when iA = 455 else
          "000111000000000"  when iA = 456 else
          "000010000000100"  when iA = 457 else
          "010110111001111"  when iA = 458 else
          "000010100100100"  when iA = 459 else
          "100000100000100"  when iA = 460 else
          "000111100100000"  when iA = 461 else
          "010000111001111"  when iA = 462 else
          "000010000000000"  when iA = 463 else
          "100000000000000"  when iA = 464 else
          "110000000011000"  when iA = 465 else
          "000110000000000"  when iA = 466 else
          "110000000100000"  when iA = 467 else
          "000010000000000"  when iA = 468 else
          "100000000000000"  when iA = 469 else
          "000000011000000"  when iA = 470 else
          "001000001000000"  when iA = 471 else
          "001000001001000"  when iA = 472 else
          "001000001001000"  when iA = 473 else
          "000110001001000"  when iA = 474 else
          "000110000000000"  when iA = 475 else
          "000110000000000"  when iA = 476 else
          "100000010000000"  when iA = 477 else
          "010010111100110"  when iA = 478 else
          "000010100010011"  when iA = 479 else
          "010001111100100"  when iA = 480 else
          "000001010000001"  when iA = 481 else
          "100000010000010"  when iA = 482 else
          "010001010101011"  when iA = 483 else
          "000110000000000"  when iA = 484 else
          "010000111011101"  when iA = 485 else
          "000000010010000"  when iA = 486 else
          "010110010101011"  when iA = 487 else
          "010000000000000"  when iA = 488 else
          "010000010101011"  when iA = 489 else
          "000010000000000"  when iA = 490 else
          "000010000000000"  when iA = 491 else
          "000010001001001"  when iA = 492 else
          "000010010010010"  when iA = 493 else
          "000010011011011"  when iA = 494 else
          "000010100100100"  when iA = 495 else
          "000010110110110"  when iA = 496 else
          "010000111101011"  when iA = 497 else
          "000000000000000";
end Behavioral;
------------------------------------------------------------------
